library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity multiplexer64 is
Port (P0,P1,P2,P3,P4,P5,P6,P7,P8,P9,P10,P11,P12,P13,P14,P15,P16,P17,P18,P19,P20,P21,P22,P23,P24,P25,P26,P27,P28,P29,P30,P31,P32,P33,P34,P35,P36,P37,P38,P39,P40,P41,P42,P43,P44,P45,P46,P47,P48,P49,P50,P51,P52,P53,P54,P55,P56,P57,P58,P59,P60,P61,P62,P63: inout std_logic_vector(15 downto 0);
      EN: in std_logic;
      Port_on_Databus: in std_logic;
    Data_on_Port: in std_logic;
PortSel:in STD_LOGIC_VECTOR (5 downto 0);
  
y : out STD_LOGIC_vector(15 downto 0);
yi : in STD_LOGIC_vector(15 downto 0));
end multiplexer64;
architecture Behavioral of multiplexer64 is
begin
process (EN,Data_on_Port,Port_on_Databus,P0,P1,P2,P3,P4,P5,P6,P7,P8,P9,P10,P11,P12,P13,P14,P15,P16,P17,P18,P19,P20,P21,P22,P23,P24,P25,P26,P27,P28,P29,P30,P31,P32,P33,P34,P35,P36,P37,P38,P39,P40,P41,P42,P43,P44,P45,P46,P47,P48,P49,P50,P51,P52,P53,P54,P55,P56,P57,P58,P59,P60,P61,P62,P63,PortSel)
begin
   
 if Port_on_Databus='1'   then
  
     
case PortSel is

when "000000"=>y<=P0;
when "000001"=>y<=P1;
when "000010"=>y<=P2;
when "000011"=>y<=P3;
when "000100"=>y<=P4;
when "000101"=>y<=P5;
when "000110"=>y<=P6;
when "000111"=>y<=P7;
when "001000"=>y<=P8;
when "001001"=>y<=P9;
when "001010"=>y<=P10;
when "001011"=>y<=P11;
when "001100"=>y<=P12;
when "001101"=>y<=P13;
when "001110"=>y<=P14;
when "001111"=>y<=P15;
when "010000"=>y<=P16;
when "010001"=>y<=P17;
when "010010"=>y<=P18;
when "010011"=>y<=P19;
when "010100"=>y<=P20;
when "010101"=>y<=P21;
when "010110"=>y<=P22;
when "010111"=>y<=P23;
when "011000"=>y<=P24;
when "011001"=>y<=P25;
when "011010"=>y<=P26;
when "011011"=>y<=P27;
when "011100"=>y<=P28;
when "011101"=>y<=P29;
when "011110"=>y<=P30;
when "011111"=>y<=P31;
when "100000"=>y<=P32;
when "100001"=>y<=P33;
when "100010"=>y<=P34;
when "100011"=>y<=P35;
when "100100"=>y<=P36;
when "100101"=>y<=P37;
when "100110"=>y<=P38;
when "100111"=>y<=P39;
when "101000"=>y<=P40;
when "101001"=>y<=P41;
when "101010"=>y<=P42;
when "101011"=>y<=P43;
when "101100"=>y<=P44;
when "101101"=>y<=P45;
when "101110"=>y<=P46;
when "101111"=>y<=P47;
when "110000"=>y<=P48;
when "110001"=>y<=P49;
when "110010"=>y<=P50;
when "110011"=>y<=P51;
when "110100"=>y<=P52;
when "110101"=>y<=P53;
when "110110"=>y<=P54;
when "110111"=>y<=P55;
when "111000"=>y<=P56;
when "111001"=>y<=P57;
when "111010"=>y<=P58;
when "111011"=>y<=P59;
when "111100"=>y<=P60;
when "111101"=>y<=P61;
when "111110"=>y<=P62;
when "111111"=>y<=P63;   
when others=> null;
end case;
else 
if Data_on_Port='1' and EN='1'  then
  case PortSel is
when "000000"=> P0<= yi;
when "000001"=> P1<= yi;
when "000010"=> P2<= yi;
when "000011"=> P3<= yi;
when "000100"=> P4<= yi;
when "000101"=> P5<= yi;
when "000110"=> P6<= yi;
when "000111"=> P7<= yi;
when "001000"=> P8<= yi;
when "001001"=> P9<= yi;
when "001010"=> P10<= yi;
when "001011"=> P11<= yi;
when "001100"=> P12<= yi;
when "001101"=> P13<= yi;
when "001110"=> P14<= yi;
when "001111"=> P15<= yi;
when "010000"=> P16<= yi;
when "010001"=> P17<= yi;
when "010010"=> P18<= yi;
when "010011"=> P19<= yi;
when "010100"=> P20<= yi;
when "010101"=> P21<= yi;
when "010110"=> P22<= yi;
when "010111"=> P23<= yi;
when "011000"=> P24<= yi;
when "011001"=> P25<= yi;
when "011010"=> P26<= yi;
when "011011"=> P27<= yi;
when "011100"=> P28<= yi;
when "011101"=> P29<= yi;
when "011110"=> P30<= yi;
when "011111"=> P31<= yi;
when "100000"=> P32<= yi;
when "100001"=> P33<= yi;
when "100010"=> P34<= yi;
when "100011"=> P35<= yi;
when "100100"=> P36<= yi;
when "100101"=> P37<= yi;
when "100110"=> P38<= yi;
when "100111"=> P39<= yi;
when "101000"=> P40<= yi;
when "101001"=> P41<= yi;
when "101010"=> P42<= yi;
when "101011"=> P43<= yi;
when "101100"=> P44<= yi;
when "101101"=> P45<= yi;
when "101110"=> P46<= yi;
when "101111"=> P47<= yi;
when "110000"=> P48<= yi;
when "110001"=> P49<= yi;
when "110010"=> P50<= yi;
when "110011"=> P51<= yi;
when "110100"=> P52<= yi;
when "110101"=> P53<= yi;
when "110110"=> P54<= yi;
when "110111"=> P55<= yi;
when "111000"=> P56<= yi;
when "111001"=> P57<= yi;
when "111010"=> P58<= yi;
when "111011"=> P59<= yi;
when "111100"=> P60<= yi;
when "111101"=> P61<= yi;
when "111110"=> P62<= yi;
when "111111"=> P63<= yi;
  when others=> null;
end case;
  
else
  case PortSel is
when "000000"=> P0<= (others => 'Z');
when "000001"=> P1<= (others => 'Z');
when "000010"=> P2<= (others => 'Z');
when "000011"=> P3<= (others => 'Z');
when "000100"=> P4<= (others => 'Z');
when "000101"=> P5<= (others => 'Z');
when "000110"=> P6<= (others => 'Z');
when "000111"=> P7<= (others => 'Z');
when "001000"=> P8<= (others => 'Z');
when "001001"=> P9<= (others => 'Z');
when "001010"=> P10<= (others => 'Z');
when "001011"=> P11<= (others => 'Z');
when "001100"=> P12<= (others => 'Z');
when "001101"=> P13<= (others => 'Z');
when "001110"=> P14<= (others => 'Z');
when "001111"=> P15<= (others => 'Z');
when "010000"=> P16<= (others => 'Z');
when "010001"=> P17<= (others => 'Z');
when "010010"=> P18<= (others => 'Z');
when "010011"=> P19<= (others => 'Z');
when "010100"=> P20<= (others => 'Z');
when "010101"=> P21<= (others => 'Z');
when "010110"=> P22<= (others => 'Z');
when "010111"=> P23<= (others => 'Z');
when "011000"=> P24<= (others => 'Z');
when "011001"=> P25<= (others => 'Z');
when "011010"=> P26<= (others => 'Z');
when "011011"=> P27<= (others => 'Z');
when "011100"=> P28<= (others => 'Z');
when "011101"=> P29<= (others => 'Z');
when "011110"=> P30<= (others => 'Z');
when "011111"=> P31<= (others => 'Z');
when "100000"=> P32<= (others => 'Z');
when "100001"=> P33<= (others => 'Z');
when "100010"=> P34<= (others => 'Z');
when "100011"=> P35<= (others => 'Z');
when "100100"=> P36<= (others => 'Z');
when "100101"=> P37<= (others => 'Z');
when "100110"=> P38<= (others => 'Z');
when "100111"=> P39<= (others => 'Z');
when "101000"=> P40<= (others => 'Z');
when "101001"=> P41<= (others => 'Z');
when "101010"=> P42<= (others => 'Z');
when "101011"=> P43<= (others => 'Z');
when "101100"=> P44<= (others => 'Z');
when "101101"=> P45<= (others => 'Z');
when "101110"=> P46<= (others => 'Z');
when "101111"=> P47<= (others => 'Z');
when "110000"=> P48<= (others => 'Z');
when "110001"=> P49<= (others => 'Z');
when "110010"=> P50<= (others => 'Z');
when "110011"=> P51<= (others => 'Z');
when "110100"=> P52<= (others => 'Z');
when "110101"=> P53<= (others => 'Z');
when "110110"=> P54<= (others => 'Z');
when "110111"=> P55<= (others => 'Z');
when "111000"=> P56<= (others => 'Z');
when "111001"=> P57<= (others => 'Z');
when "111010"=> P58<= (others => 'Z');
when "111011"=> P59<= (others => 'Z');
when "111100"=> P60<= (others => 'Z');
when "111101"=> P61<= (others => 'Z');
when "111110"=> P62<= (others => 'Z');
when "111111"=> P63<= (others => 'Z');
  when others=> null;
end case;
  end if;
end if;
end process;
End Behavioral;