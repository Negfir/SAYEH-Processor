library IEEE;
use IEEE.std_logic_1164.ALL;
ENTITY Main_TB is
END Main_TB;
ARCHITECTURE simulate OF Main_TB IS
  
COMPONENT Main IS
	PORT (P0,P1,P2,P3,P4,P5,P6,P7,P8,P9,P10,P11,P12,P13,P14,P15,P16,P17,P18,P19,P20,P21,P22,P23,P24,P25,P26,P27,P28,P29,P30,P31,P32,P33,P34,P35,P36,P37,P38,P39,P40,P41,P42,P43,P44,P45,P46,P47,P48,P49,P50,P51,P52,P53,P54,P55,P56,P57,P58,P59,P60,P61,P62,P63 : inout std_logic_vector(15 downto 0);
  External_Reset : in std_logic;
	clk: in std_logic);
	
	  end COMPONENT;  

signal clk, reset : std_logic := '0';
signal P0,P1,P2,P3,P4,P5,P6,P7,P8,P9,P10,P11,P12,P13,P14,P15,P16,P17,P18,P19,P20,P21,P22,P23,P24,P25,P26,P27,P28,P29,P30,P31,P32,P33,P34,P35,P36,P37,P38,P39,P40,P41,P42,P43,P44,P45,P46,P47,P48,P49,P50,P51,P52,P53,P54,P55,P56,P57,P58,P59,P60,P61,P62,P63 :  std_logic_vector(15 downto 0):="0000000000000000";

BEGIN

Sayeh : main port map (P0,P1,P2,P3,P4,P5,P6,P7,P8,P9,P10,P11,P12,P13,P14,P15,P16,P17,P18,P19,P20,P21,P22,P23,P24,P25,P26,P27,P28,P29,P30,P31,P32,P33,P34,P35,P36,P37,P38,P39,P40,P41,P42,P43,P44,P45,P46,P47,P48,P49,P50,P51,P52,P53,P54,P55,P56,P57,P58,P59,P60,P61,P62,P63, reset, clk);
	p16<="0011011100011111";
	reset <= '1', '0' after 10 ns;
	clk <= not clk after 50 ns;
	
END simulate;